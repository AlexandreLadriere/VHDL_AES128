------------------------------------------------------------------------------------------------
-- Author:			Alexandre LADRIERE
-- Name:			InvSubBytes.vhd
-- Date of creation:		14/11/2018
-- Date of modification:	14/11/2018
-- Description:			Test bench for th inversion of the ShiftRows function
------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
library AESLibrary;
use AESLibrary.state_definition_package.all;
library source;

entity InvShiftRows_tb is 
end entity InvShiftRows_tb;

architecture InvShiftRows_tb_arch of InvShiftRows_tb is
	component InvShiftRows
		port (
			invshiftrows_i : in type_state; -- matrice d'entree
			invshiftrows_o : out type_state -- matrice de sortie
		);
	end component;
	
	signal invshiftrows_is : type_state := ((x"06",x"85",x"a6",x"61"),(x"fb",x"06",x"54",x"09"),(x"5f",x"ca",x"99",x"c1"),(x"74",x"5b",x"8e",x"56"));
	signal invshiftrows_os : type_state;
	
	begin
	-- Device Under Test
	DUT : InvShiftRows
		port map (
			invshiftrows_i => invshiftrows_is,
			invshiftrows_o => invshiftrows_os
		);
end architecture InvShiftRows_tb_arch;

configuration InvShiftRows_tb_conf of InvShiftRows_tb is
	for InvShiftRows_tb_arch
		for DUT : InvShiftRows
			use entity source.InvShiftRows(InvShiftRows_arch);
		end for;
	end for;
end InvShiftRows_tb_conf;
